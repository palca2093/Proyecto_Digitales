module byte_striping();
















endmodule
